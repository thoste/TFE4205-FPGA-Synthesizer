
module clocks (
	clk_0_clk,
	reset_0_reset_n,
	reset_1_reset_n,
	clk_1_clk,
	clock_27_clk_clk,
	clock_27_reset_reset_n,
	clock_25_clk,
	clock_25_reset_reset_n);	

	input		clk_0_clk;
	input		reset_0_reset_n;
	input		reset_1_reset_n;
	input		clk_1_clk;
	output		clock_27_clk_clk;
	output		clock_27_reset_reset_n;
	output		clock_25_clk;
	output		clock_25_reset_reset_n;
endmodule
