// clocks.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module clocks (
		input  wire  clk_0_clk,              //          clk_0.clk
		input  wire  clk_1_clk,              //          clk_1.clk
		output wire  clock_25_clk,           //       clock_25.clk
		output wire  clock_25_reset_reset_n, // clock_25_reset.reset_n
		output wire  clock_27_clk_clk,       //   clock_27_clk.clk
		output wire  clock_27_reset_reset_n, // clock_27_reset.reset_n
		input  wire  reset_0_reset_n,        //        reset_0.reset_n
		input  wire  reset_1_reset_n         //        reset_1.reset_n
	);

	assign clock_27_clk_clk = clk_0_clk;

	assign clock_25_clk = clk_1_clk;

	assign clock_27_reset_reset_n = reset_0_reset_n;

	assign clock_25_reset_reset_n = reset_1_reset_n;

endmodule
